/*                                                                      
 Copyright 2025 Yusen Wang @yusen.w@qq.com
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
 Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */

`include "defines.v"

// 将译码结果向执行模块传递
module id_ex (

    input wire                        clk,
    input wire                        rst,
    // 输入
    input wire [                31:0] inst_i,          // 指令内容
    input wire [`INST_ADDR_WIDTH-1:0] inst_addr_i,     // 指令地址
    input wire                        reg_we_i,        // 写通用寄存器标志
    input wire [ `REG_ADDR_WIDTH-1:0] reg_waddr_i,     // 写通用寄存器地址
    input wire [ `REG_DATA_WIDTH-1:0] reg1_rdata_i,    // 通用寄存器1读数据
    input wire [ `REG_DATA_WIDTH-1:0] reg2_rdata_i,    // 通用寄存器2读数据
    input wire                        csr_we_i,        // 写CSR寄存器标志
    input wire [ `BUS_ADDR_WIDTH-1:0] csr_waddr_i,     // 写CSR寄存器地址
    input wire [ `REG_DATA_WIDTH-1:0] csr_rdata_i,     // CSR寄存器读数据
    input wire [  `DECINFO_WIDTH-1:0] dec_info_bus_i,
    input wire [                31:0] dec_imm_i,

    input wire [`Hold_Flag_Bus] hold_flag_i,  // 流水线暂停标志

    output wire [`INST_DATA_WIDTH-1:0] inst_o,         // 指令内容
    output wire [`INST_ADDR_WIDTH-1:0] inst_addr_o,    // 指令地址
    output wire                        reg_we_o,       // 写通用寄存器标志
    output wire [ `REG_ADDR_WIDTH-1:0] reg_waddr_o,    // 写通用寄存器地址
    output wire [ `REG_DATA_WIDTH-1:0] reg1_rdata_o,   // 通用寄存器1读数据
    output wire [ `REG_DATA_WIDTH-1:0] reg2_rdata_o,   // 通用寄存器2读数据
    output wire                        csr_we_o,       // 写CSR寄存器标志
    output wire [ `REG_DATA_WIDTH-1:0] csr_rdata_o,    // CSR寄存器读数据
    output wire [                31:0] dec_imm_o,      // 立即数
    output wire [ `BUS_ADDR_WIDTH-1:0] csr_waddr_o,    // 写CSR寄存器地址
    output wire [  `DECINFO_WIDTH-1:0] dec_info_bus_o  // 译码信息总线
);

    wire                        hold_en = (hold_flag_i >= `Hold_Id);

    wire [`INST_DATA_WIDTH-1:0] inst;
    gen_pipe_dff #(32) inst_ff (
        clk,
        rst,
        hold_en,
        `INST_NOP,
        inst_i,
        inst
    );
    assign inst_o = inst;

    wire [`INST_ADDR_WIDTH-1:0] inst_addr;
    gen_pipe_dff #(32) inst_addr_ff (
        clk,
        rst,
        hold_en,
        `ZeroWord,
        inst_addr_i,
        inst_addr
    );
    assign inst_addr_o = inst_addr;

    wire reg_we;
    gen_pipe_dff #(1) reg_we_ff (
        clk,
        rst,
        hold_en,
        `WriteDisable,
        reg_we_i,
        reg_we
    );
    assign reg_we_o = reg_we;

    wire [`REG_ADDR_WIDTH-1:0] reg_waddr;
    gen_pipe_dff #(5) reg_waddr_ff (
        clk,
        rst,
        hold_en,
        `ZeroReg,
        reg_waddr_i,
        reg_waddr
    );
    assign reg_waddr_o = reg_waddr;

    wire [`REG_DATA_WIDTH-1:0] reg1_rdata;
    gen_pipe_dff #(32) reg1_rdata_ff (
        clk,
        rst,
        hold_en,
        `ZeroWord,
        reg1_rdata_i,
        reg1_rdata
    );
    assign reg1_rdata_o = reg1_rdata;

    wire [`REG_DATA_WIDTH-1:0] reg2_rdata;
    gen_pipe_dff #(32) reg2_rdata_ff (
        clk,
        rst,
        hold_en,
        `ZeroWord,
        reg2_rdata_i,
        reg2_rdata
    );
    assign reg2_rdata_o = reg2_rdata;

    wire csr_we;
    gen_pipe_dff #(1) csr_we_ff (
        clk,
        rst,
        hold_en,
        `WriteDisable,
        csr_we_i,
        csr_we
    );
    assign csr_we_o = csr_we;

    wire [`BUS_ADDR_WIDTH-1:0] csr_waddr;
    gen_pipe_dff #(32) csr_waddr_ff (
        clk,
        rst,
        hold_en,
        `ZeroWord,
        csr_waddr_i,
        csr_waddr
    );
    assign csr_waddr_o = csr_waddr;

    wire [`REG_DATA_WIDTH-1:0] csr_rdata;
    gen_pipe_dff #(32) csr_rdata_ff (
        clk,
        rst,
        hold_en,
        `ZeroWord,
        csr_rdata_i,
        csr_rdata
    );
    assign csr_rdata_o = csr_rdata;

    // 新增译码信息总线传递
    wire [`DECINFO_WIDTH-1:0] dec_info_bus;
    gen_pipe_dff #(`DECINFO_WIDTH) dec_info_bus_ff (
        clk,
        rst,
        hold_en,
        `ZeroWord,
        dec_info_bus_i,
        dec_info_bus
    );
    assign dec_info_bus_o = dec_info_bus;

    // 新增立即数传递
    wire [31:0] dec_imm;
    gen_pipe_dff #(32) dec_imm_ff (
        clk,
        rst,
        hold_en,
        `ZeroWord,
        dec_imm_i,
        dec_imm
    );
    assign dec_imm_o = dec_imm;

endmodule
