/*                                                                      
 Copyright 2025 Yusen Wang @yusen.w@qq.com
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
 Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */

`include "defines.svh"

// 控制模块
// 发出跳转、暂停流水线信号
module ctrl (

    input wire rst_n,

    // from ex
    input wire                        jump_flag_i,
    input wire [`INST_ADDR_WIDTH-1:0] jump_addr_i,
    input wire                        hold_flag_ex_i,

    // from mems arbiter
    input wire hold_flag_mems_i,

    // from clint
    input wire hold_flag_clint_i,

    // from HDU - 新增
    input wire hold_flag_hdu_i,

    output reg [`Hold_Flag_Bus] hold_flag_o,

    // to pc_reg
    output reg                        jump_flag_o,
    output reg [`INST_ADDR_WIDTH-1:0] jump_addr_o

);


    always @(*) begin
        jump_addr_o = jump_addr_i;
        jump_flag_o = jump_flag_i;
        // 默认不暂停
        hold_flag_o = `Hold_None;
        // 按优先级处理不同模块的请求
        if (jump_flag_i == `JumpEnable || hold_flag_ex_i == `HoldEnable || 
            hold_flag_clint_i == `HoldEnable) begin  // 新增HDU暂停条件
            // 暂停整条流水线
            hold_flag_o = `Hold_Id;
        end else if (hold_flag_mems_i == `HoldEnable || hold_flag_hdu_i == `HoldEnable) begin
            // 暂停PC，即取指地址不变
            hold_flag_o = `Hold_Pc;
        end else begin
            hold_flag_o = `Hold_None;
        end
    end

endmodule
