/*         
 The MIT License (MIT)

 Copyright © 2025 Yusen Wang @yusen.w@qq.com
                                                                         
 Permission is hereby granted, free of charge, to any person obtaining a copy
 of this software and associated documentation files (the "Software"), to deal
 in the Software without restriction, including without limitation the rights
 to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 copies of the Software, and to permit persons to whom the Software is
 furnished to do so, subject to the following conditions:
                                                                         
 The above copyright notice and this permission notice shall be included in all
 copies or substantial portions of the Software.
                                                                         
 THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 SOFTWARE.
 */

`include "defines.svh"

// 冒险检测单元 - 处理长指令的RAW和WAW相关性
module hdu (
    input wire clk,   // 时钟
    input wire rst_n, // 复位信号，低电平有效

    // 新指令信息
    input wire                          inst_valid,  // 新长指令有效
    input wire [   `REG_ADDR_WIDTH-1:0] rd_addr,     // 新指令写寄存器地址
    input wire [   `REG_ADDR_WIDTH-1:0] rs1_addr,    // 新指令读寄存器1地址
    input wire [   `REG_ADDR_WIDTH-1:0] rs2_addr,    // 新指令读寄存器2地址
    input wire                          rd_we,       // 新指令是否写寄存器
    input wire                          rs1_re,      // 是否检测rs1
    input wire                          rs2_re,      // 是否检测rs2
    input wire [`EX_INFO_BUS_WIDTH-1:0] ex_info_bus, // 新增：指令ex单元类型

    // 长指令完成信号
    input wire                        commit_valid_i,  // 长指令执行完成有效信号
    input wire [`COMMIT_ID_WIDTH-1:0] commit_id_i,     // 执行完成的长指令ID

    // 控制信号
    output wire hazard_stall_o,  // 暂停流水线信号
    output wire [`COMMIT_ID_WIDTH-1:0] commit_id_o,  // 为新的长指令分配的ID
    output wire long_inst_atom_lock_o,  // 原子锁信号，FIFO中有未销毁的长指令时为1
    output wire alu_pass_op1_o,  // ALU rs1 RAW冒险旁路前递，特判放行
    output wire alu_pass_op2_o,  // ALU rs2 RAW冒险旁路前递，特判放行
    output wire mul_pass_op1_o,  // MUL rs1 RAW冒险旁路前递
    output wire mul_pass_op2_o,  // MUL rs2 RAW冒险旁路前递
    output wire div_pass_op1_o,  // DIV rs1 RAW冒险旁路前递
    output wire div_pass_op2_o,  // DIV rs2 RAW冒险旁路前递
    output wire csr_pass_op1_o  // CSR rs1 RAW冒险旁路前递
);

    // 定义FIFO表项结构
    typedef struct packed {
        logic [`REG_ADDR_WIDTH-1:0] rd_addr;
        logic [`EX_INFO_BUS_WIDTH-1:0] exu_type;
    } fifo_entry_t;

    reg [7:0] fifo_valid;  // 有效位，深度8
    fifo_entry_t fifo_entry[0:7];  // 存储表项结构体，深度8

    // 冒险检测信号
    reg raw_hazard;  // 读后写冒险
    reg waw_hazard;  // 写后写冒险
    wire hazard;  // 总冒险信号

    // ALU RAW冒险掩码及其对应ID
    reg [7:0] alu_raw_mask;
    reg [2:0] alu_raw_mask_id;  // 记录当前mask对应的commit_id

    // RAW冒险对象指示
    reg alu_raw_rs1, alu_raw_rs2;
    reg mul_raw_rs1, mul_raw_rs2;
    reg div_raw_rs1, div_raw_rs2;
    reg        csr_raw_rs1;

    // RAW冒险向量
    wire [7:0] raw_hazard_vec;
    wire [7:0] waw_hazard_vec;
    wire [7:0] masked_raw_hazard_vec;

    wire       is_alu_inst = (ex_info_bus == `EX_INFO_ALU);
    wire       is_mul_inst = (ex_info_bus == `EX_INFO_MUL);
    wire       is_div_inst = (ex_info_bus == `EX_INFO_DIV);
    wire       is_csr_inst = (ex_info_bus == `EX_INFO_CSR);
    wire       is_alu_bypass_inst = (ex_info_bus[`EX_INFO_BYPASS_BIT] == 1'b0);

    genvar i;
    generate
        for (i = 0; i < 8; i = i + 1) begin : hazard_vec_gen
            assign raw_hazard_vec[i] = fifo_valid[i] && !(commit_valid_i && commit_id_i == i) &&
                ((rs1_re && rs1_addr == fifo_entry[i].rd_addr) || (rs2_re && rs2_addr == fifo_entry[i].rd_addr));
            // waw检测：只有exu_type不同才算冲突
            assign waw_hazard_vec[i] = fifo_valid[i] && !(commit_valid_i && commit_id_i == i) &&
                (rd_we && rd_addr == fifo_entry[i].rd_addr && ex_info_bus != fifo_entry[i].exu_type);
        end
    endgenerate

    // RAW冒险掩码更新
    always @(posedge clk or negedge rst_n) begin
        if (~rst_n) begin
            alu_raw_mask    <= 8'hFF;
            alu_raw_mask_id <= 3'd0;
        end else begin
            // 清除已完成的长指令
            if (commit_valid_i && (alu_raw_mask_id == commit_id_i)) begin
                alu_raw_mask    <= 8'hFF;
                alu_raw_mask_id <= 3'd0;
            end
            // 添加新的ALU写寄存器指令，分配mask并记录id
            if (inst_valid && ~hazard && is_alu_inst && rd_we) begin
                alu_raw_mask    <= ~(8'b1 << commit_id_o);
                alu_raw_mask_id <= commit_id_o;
            end
        end
    end

    assign masked_raw_hazard_vec = is_alu_bypass_inst ? (raw_hazard_vec & alu_raw_mask) : raw_hazard_vec;
    // RAW冒险输出（掩码屏蔽新分配ID）
    assign raw_hazard = |masked_raw_hazard_vec;
    assign waw_hazard = |waw_hazard_vec;

    // 只有在有新指令且存在冒险时才暂停流水线
    assign hazard = (raw_hazard || waw_hazard);
    assign hazard_stall_o = hazard || (&fifo_valid);  // 如果FIFO已满也暂停流水线

    // 为新的长指令分配ID - 使用assign语句
    assign commit_id_o = (inst_valid && ~hazard) ?
        ( ~fifo_valid[0] ? 0 :
          ~fifo_valid[1] ? 1 :
          ~fifo_valid[2] ? 2 :
          ~fifo_valid[3] ? 3 :
          ~fifo_valid[4] ? 4 :
          ~fifo_valid[5] ? 5 :
          ~fifo_valid[6] ? 6 :
          ~fifo_valid[7] ? 7 : 0 ) : 0;

    // 更新FIFO
    always @(posedge clk or negedge rst_n) begin
        if (~rst_n) begin
            // 复位时清空FIFO
            for (int i = 0; i < 8; i = i + 1) begin
                fifo_valid[i]          <= 1'b0;
                fifo_entry[i].rd_addr  <= 5'h0;
                fifo_entry[i].exu_type <= {`EX_INFO_BUS_WIDTH{1'b0}};
            end
        end else begin
            // 清除已完成的长指令
            if (commit_valid_i) begin
                fifo_valid[commit_id_i] <= 1'b0;
            end

            // 添加新的长指令到FIFO
            if (inst_valid && ~hazard) begin
                fifo_valid[commit_id_o]          <= 1'b1;
                fifo_entry[commit_id_o].rd_addr  <= rd_addr;
                fifo_entry[commit_id_o].exu_type <= ex_info_bus;
            end
        end
    end

    // RAW冒险对象检测（对ALU/MUL/DIV/CSR指令有效）
    always @(*) begin
        alu_raw_rs1 = 1'b0;
        alu_raw_rs2 = 1'b0;
        mul_raw_rs1 = 1'b0;
        mul_raw_rs2 = 1'b0;
        div_raw_rs1 = 1'b0;
        div_raw_rs2 = 1'b0;
        csr_raw_rs1 = 1'b0;
        if (is_alu_inst) begin
            // 只需检查alu_raw_mask_id对应的FIFO表项，且只关心通道一写回
            if (fifo_valid[alu_raw_mask_id] && alu_raw_mask != 8'hFF &&
                !(commit_valid_i && commit_id_i == alu_raw_mask_id)) begin
                if (rs1_re && rs1_addr == fifo_entry[alu_raw_mask_id].rd_addr) alu_raw_rs1 = 1'b1;
                if (rs2_re && rs2_addr == fifo_entry[alu_raw_mask_id].rd_addr) alu_raw_rs2 = 1'b1;
            end
        end
        if (is_mul_inst) begin
            if (fifo_valid[alu_raw_mask_id] && alu_raw_mask != 8'hFF &&
                !(commit_valid_i && commit_id_i == alu_raw_mask_id)) begin
                if (rs1_re && rs1_addr == fifo_entry[alu_raw_mask_id].rd_addr) mul_raw_rs1 = 1'b1;
                if (rs2_re && rs2_addr == fifo_entry[alu_raw_mask_id].rd_addr) mul_raw_rs2 = 1'b1;
            end
        end
        if (is_div_inst) begin
            if (fifo_valid[alu_raw_mask_id] && alu_raw_mask != 8'hFF &&
                !(commit_valid_i && commit_id_i == alu_raw_mask_id)) begin
                if (rs1_re && rs1_addr == fifo_entry[alu_raw_mask_id].rd_addr) div_raw_rs1 = 1'b1;
                if (rs2_re && rs2_addr == fifo_entry[alu_raw_mask_id].rd_addr) div_raw_rs2 = 1'b1;
            end
        end
        if (is_csr_inst) begin
            if (fifo_valid[alu_raw_mask_id] && alu_raw_mask != 8'hFF &&
                !(commit_valid_i && commit_id_i == alu_raw_mask_id)) begin
                if (rs1_re && rs1_addr == fifo_entry[alu_raw_mask_id].rd_addr) csr_raw_rs1 = 1'b1;
            end
        end
    end

    assign alu_pass_op1_o        = alu_raw_rs1;
    assign alu_pass_op2_o        = alu_raw_rs2;
    assign mul_pass_op1_o        = mul_raw_rs1;
    assign mul_pass_op2_o        = mul_raw_rs2;
    assign div_pass_op1_o        = div_raw_rs1;
    assign div_pass_op2_o        = div_raw_rs2;
    assign csr_pass_op1_o        = csr_raw_rs1;

    // 生成原子锁信号 - 当FIFO中有任何一个有效的长指令时为1
    assign long_inst_atom_lock_o = |fifo_valid;
endmodule
