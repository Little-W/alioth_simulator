/*
 The MIT License (MIT)

 Copyright © 2025 Yusen Wang @yusen.w@qq.com
                                                                         
 Permission is hereby granted, free of charge, to any person obtaining a copy
 of this software and associated documentation files (the "Software"), to deal
 in the Software without restriction, including without limitation the rights
 to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 copies of the Software, and to permit persons to whom the Software is
 furnished to do so, subject to the following conditions:
                                                                         
 The above copyright notice and this permission notice shall be included in all
 copies or substantial portions of the Software.
                                                                         
 THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 SOFTWARE.
 */

`include "defines.svh"

module axi_interconnect #(
    parameter int IMEM_ADDR_WIDTH = 16,
    parameter int DMEM_ADDR_WIDTH = 16,
    parameter int DATA_WIDTH      = 32,
    parameter int C_AXI_ID_WIDTH   = 2,
    parameter int C_AXI_DATA_WIDTH = 32,
    parameter int C_AXI_ADDR_WIDTH = 32,
    parameter int C_OM0_AXI_ADDR_WIDTH = 32,
    parameter int C_OM0_AXI_DATA_WIDTH = 32,
    parameter int C_OM1_AXI_ADDR_WIDTH = 32,
    parameter int C_OM1_AXI_DATA_WIDTH = 32,
    parameter int C_OM2_AXI_ADDR_WIDTH = 32,
    parameter int C_OM2_AXI_DATA_WIDTH = 32
) (
    // 全局信号
    input wire clk,
    input wire rst_n,

    // Master 0 接口
    input  wire [C_AXI_ID_WIDTH-1:0]     M0_AXI_ARID,
    input  wire [C_AXI_ADDR_WIDTH-1:0]  M0_AXI_ARADDR,
    input  wire [7:0]                    M0_AXI_ARLEN,
    input  wire [2:0]                    M0_AXI_ARSIZE,
    input  wire [1:0]                    M0_AXI_ARBURST,
    input  wire                          M0_AXI_ARLOCK,
    input  wire [3:0]                    M0_AXI_ARCACHE,
    input  wire [2:0]                    M0_AXI_ARPROT,
    input  wire [3:0]                    M0_AXI_ARQOS,
    input  wire [3:0]                    M0_AXI_ARUSER,
    input  wire                          M0_AXI_ARVALID,
    output wire                          M0_AXI_ARREADY,
    output wire [C_AXI_ID_WIDTH-1:0]     M0_AXI_RID,
    output wire [C_AXI_DATA_WIDTH-1:0]  M0_AXI_RDATA,
    output wire [1:0]                    M0_AXI_RRESP,
    output wire                          M0_AXI_RLAST,
    output wire [3:0]                    M0_AXI_RUSER,
    output wire                          M0_AXI_RVALID,
    input  wire                          M0_AXI_RREADY,

    // Master 1 接口
    input  wire [C_AXI_ID_WIDTH-1:0]     M1_AXI_AWID,
    input  wire [C_AXI_ADDR_WIDTH-1:0]  M1_AXI_AWADDR,
    input  wire [7:0]                    M1_AXI_AWLEN,
    input  wire [2:0]                    M1_AXI_AWSIZE,
    input  wire [1:0]                    M1_AXI_AWBURST,
    input  wire                          M1_AXI_AWLOCK,
    input  wire [3:0]                    M1_AXI_AWCACHE,
    input  wire [2:0]                    M1_AXI_AWPROT,
    input  wire [3:0]                    M1_AXI_AWQOS,
    input  wire [3:0]                    M1_AXI_AWUSER,
    input  wire                          M1_AXI_AWVALID,
    output wire                          M1_AXI_AWREADY,
    input  wire [C_AXI_DATA_WIDTH-1:0]  M1_AXI_WDATA,
    input  wire [(C_AXI_DATA_WIDTH/8)-1:0] M1_AXI_WSTRB,
    input  wire                          M1_AXI_WLAST,
    input  wire                          M1_AXI_WVALID,
    output wire                          M1_AXI_WREADY,
    output wire [C_AXI_ID_WIDTH-1:0]     M1_AXI_BID,
    output wire [1:0]                    M1_AXI_BRESP,
    output wire                          M1_AXI_BVALID,
    input  wire                          M1_AXI_BREADY,
    input  wire [C_AXI_ID_WIDTH-1:0]     M1_AXI_ARID,
    input  wire [C_AXI_ADDR_WIDTH-1:0]  M1_AXI_ARADDR,
    input  wire [7:0]                    M1_AXI_ARLEN,
    input  wire [2:0]                    M1_AXI_ARSIZE,
    input  wire [1:0]                    M1_AXI_ARBURST,
    input  wire                          M1_AXI_ARLOCK,
    input  wire [3:0]                    M1_AXI_ARCACHE,
    input  wire [2:0]                    M1_AXI_ARPROT,
    input  wire [3:0]                    M1_AXI_ARQOS,
    input  wire [3:0]                    M1_AXI_ARUSER,
    input  wire                          M1_AXI_ARVALID,
    output wire                          M1_AXI_ARREADY,
    output wire [C_AXI_ID_WIDTH-1:0]     M1_AXI_RID,
    output wire [C_AXI_DATA_WIDTH-1:0]  M1_AXI_RDATA,
    output wire [1:0]                    M1_AXI_RRESP,
    output wire                          M1_AXI_RLAST,
    output wire [3:0]                    M1_AXI_RUSER,
    output wire                          M1_AXI_RVALID,
    input  wire                          M1_AXI_RREADY,

    // Slave 接口...
    // APB AXI-lite 接口
    output wire                                  OM0_AXI_ACLK,
    output wire                                  OM0_AXI_ARESETN,
    output wire [    C_OM0_AXI_ADDR_WIDTH-1 : 0] OM0_AXI_AWADDR,
    output wire [                         2 : 0] OM0_AXI_AWPROT,
    output wire                                  OM0_AXI_AWVALID,
    input  wire                                  OM0_AXI_AWREADY,
    output wire [    C_OM0_AXI_DATA_WIDTH-1 : 0] OM0_AXI_WDATA,
    output wire [(C_OM0_AXI_DATA_WIDTH/8)-1 : 0] OM0_AXI_WSTRB,
    output wire                                  OM0_AXI_WVALID,
    input  wire                                  OM0_AXI_WREADY,
    input  wire [                         1 : 0] OM0_AXI_BRESP,
    input  wire                                  OM0_AXI_BVALID,
    output wire                                  OM0_AXI_BREADY,
    output wire [    C_OM0_AXI_ADDR_WIDTH-1 : 0] OM0_AXI_ARADDR,
    output wire [                         2 : 0] OM0_AXI_ARPROT,
    output wire                                  OM0_AXI_ARVALID,
    input  wire                                  OM0_AXI_ARREADY,
    input  wire [    C_OM0_AXI_DATA_WIDTH-1 : 0] OM0_AXI_RDATA,
    input  wire [                         1 : 0] OM0_AXI_RRESP,
    input  wire                                  OM0_AXI_RVALID,
    output wire                                  OM0_AXI_RREADY,
    // CLINT AXI-lite 接口
    output wire                                  OM1_AXI_ACLK,
    output wire                                  OM1_AXI_ARESETN,
    output wire [    C_OM1_AXI_ADDR_WIDTH-1 : 0] OM1_AXI_AWADDR,
    output wire [                         2 : 0] OM1_AXI_AWPROT,
    output wire                                  OM1_AXI_AWVALID,
    input  wire                                  OM1_AXI_AWREADY,
    output wire [    C_OM1_AXI_DATA_WIDTH-1 : 0] OM1_AXI_WDATA,
    output wire [(C_OM1_AXI_DATA_WIDTH/8)-1 : 0] OM1_AXI_WSTRB,
    output wire                                  OM1_AXI_WVALID,
    input  wire                                  OM1_AXI_WREADY,
    input  wire [                         1 : 0] OM1_AXI_BRESP,
    input  wire                                  OM1_AXI_BVALID,
    output wire                                  OM1_AXI_BREADY,
    output wire [    C_OM1_AXI_ADDR_WIDTH-1 : 0] OM1_AXI_ARADDR,
    output wire [                         2 : 0] OM1_AXI_ARPROT,
    output wire                                  OM1_AXI_ARVALID,
    input  wire                                  OM1_AXI_ARREADY,
    input  wire [    C_OM1_AXI_DATA_WIDTH-1 : 0] OM1_AXI_RDATA,
    input  wire [                         1 : 0] OM1_AXI_RRESP,
    input  wire                                  OM1_AXI_RVALID,
    output wire                                  OM1_AXI_RREADY,

    // CLINT AXI-lite 接口
    output wire                                  OM2_AXI_ACLK,
    output wire                                  OM2_AXI_ARESETN,
    output wire [    C_OM2_AXI_ADDR_WIDTH-1 : 0] OM2_AXI_AWADDR,
    output wire [                         2 : 0] OM2_AXI_AWPROT,
    output wire                                  OM2_AXI_AWVALID,
    input  wire                                  OM2_AXI_AWREADY,
    output wire [    C_OM2_AXI_DATA_WIDTH-1 : 0] OM2_AXI_WDATA,
    output wire [(C_OM2_AXI_DATA_WIDTH/8)-1 : 0] OM2_AXI_WSTRB,
    output wire                                  OM2_AXI_WVALID,
    input  wire                                  OM2_AXI_WREADY,
    input  wire [                         1 : 0] OM2_AXI_BRESP,
    input  wire                                  OM2_AXI_BVALID,
    output wire                                  OM2_AXI_BREADY,
    output wire [    C_OM2_AXI_ADDR_WIDTH-1 : 0] OM2_AXI_ARADDR,
    output wire [                         2 : 0] OM2_AXI_ARPROT,
    output wire                                  OM2_AXI_ARVALID,
    input  wire                                  OM2_AXI_ARREADY,
    input  wire [    C_OM2_AXI_DATA_WIDTH-1 : 0] OM2_AXI_RDATA,
    input  wire [                         1 : 0] OM2_AXI_RRESP,
    input  wire                                  OM2_AXI_RVALID,
    output wire                                  OM2_AXI_RREADY,

    // IMEM AXI接口 (指令存储器)
    output wire [  C_AXI_ID_WIDTH-1:0] IMEM_AXI_AWID,
    output wire [C_AXI_ADDR_WIDTH-1:0] IMEM_AXI_AWADDR,
    output wire [                 7:0] IMEM_AXI_AWLEN,
    output wire [                 2:0] IMEM_AXI_AWSIZE,
    output wire [                 1:0] IMEM_AXI_AWBURST,
    output wire                        IMEM_AXI_AWLOCK,
    output wire [                 3:0] IMEM_AXI_AWCACHE,
    output wire [                 2:0] IMEM_AXI_AWPROT,
    output wire                        IMEM_AXI_AWVALID,
    input  wire                        IMEM_AXI_AWREADY,
    output wire [    C_AXI_DATA_WIDTH-1:0] IMEM_AXI_WDATA,
    output wire [(C_AXI_DATA_WIDTH/8)-1:0] IMEM_AXI_WSTRB,
    output wire                            IMEM_AXI_WLAST,
    output wire                            IMEM_AXI_WVALID,
    input  wire                            IMEM_AXI_WREADY,
    input  wire [C_AXI_ID_WIDTH-1:0] IMEM_AXI_BID,
    input  wire [               1:0] IMEM_AXI_BRESP,
    input  wire                      IMEM_AXI_BVALID,
    output wire                      IMEM_AXI_BREADY,
    output wire [  C_AXI_ID_WIDTH-1:0] IMEM_AXI_ARID,
    output wire [C_AXI_ADDR_WIDTH-1:0] IMEM_AXI_ARADDR,
    output wire [                 7:0] IMEM_AXI_ARLEN,
    output wire [                 2:0] IMEM_AXI_ARSIZE,
    output wire [                 1:0] IMEM_AXI_ARBURST,
    output wire                        IMEM_AXI_ARLOCK,
    output wire [                 3:0] IMEM_AXI_ARCACHE,
    output wire [                 2:0] IMEM_AXI_ARPROT,
    output wire                        IMEM_AXI_ARVALID,
    input  wire                        IMEM_AXI_ARREADY,
    input  wire [  C_AXI_ID_WIDTH-1:0] IMEM_AXI_RID,
    input  wire [C_AXI_DATA_WIDTH-1:0] IMEM_AXI_RDATA,
    input  wire [                 1:0] IMEM_AXI_RRESP,
    input  wire                        IMEM_AXI_RLAST,
    input  wire                        IMEM_AXI_RVALID,
    output wire                        IMEM_AXI_RREADY,

    // DMEM AXI接口 (数据存储器)
    output wire [  C_AXI_ID_WIDTH-1:0] DMEM_AXI_AWID,
    output wire [C_AXI_ADDR_WIDTH-1:0] DMEM_AXI_AWADDR,
    output wire [                 7:0] DMEM_AXI_AWLEN,
    output wire [                 2:0] DMEM_AXI_AWSIZE,
    output wire [                 1:0] DMEM_AXI_AWBURST,
    output wire                        DMEM_AXI_AWLOCK,
    output wire [                 3:0] DMEM_AXI_AWCACHE,
    output wire [                 2:0] DMEM_AXI_AWPROT,
    output wire                        DMEM_AXI_AWVALID,
    input  wire                        DMEM_AXI_AWREADY,
    output wire [    C_AXI_DATA_WIDTH-1:0] DMEM_AXI_WDATA,
    output wire [(C_AXI_DATA_WIDTH/8)-1:0] DMEM_AXI_WSTRB,
    output wire                            DMEM_AXI_WLAST,
    output wire                            DMEM_AXI_WVALID,
    input  wire                            DMEM_AXI_WREADY,
    input  wire [C_AXI_ID_WIDTH-1:0] DMEM_AXI_BID,
    input  wire [               1:0] DMEM_AXI_BRESP,
    input  wire                      DMEM_AXI_BVALID,
    output wire                      DMEM_AXI_BREADY,
    output wire [  C_AXI_ID_WIDTH-1:0] DMEM_AXI_ARID,
    output wire [C_AXI_ADDR_WIDTH-1:0] DMEM_AXI_ARADDR,
    output wire [                 7:0] DMEM_AXI_ARLEN,
    output wire [                 2:0] DMEM_AXI_ARSIZE,
    output wire [                 1:0] DMEM_AXI_ARBURST,
    output wire                        DMEM_AXI_ARLOCK,
    output wire [                 3:0] DMEM_AXI_ARCACHE,
    output wire [                 2:0] DMEM_AXI_ARPROT,
    output wire                        DMEM_AXI_ARVALID,
    input  wire                        DMEM_AXI_ARREADY,
    input  wire [  C_AXI_ID_WIDTH-1:0] DMEM_AXI_RID,
    input  wire [C_AXI_DATA_WIDTH-1:0] DMEM_AXI_RDATA,
    input  wire [                 1:0] DMEM_AXI_RRESP,
    input  wire                        DMEM_AXI_RLAST,
    input  wire                        DMEM_AXI_RVALID,
    output wire                        DMEM_AXI_RREADY,

    // DM AXI接口 (Debug Module)
    output wire [  C_AXI_ID_WIDTH-1:0] DM_AXI_AWID,
    output wire [C_AXI_ADDR_WIDTH-1:0] DM_AXI_AWADDR,
    output wire [                 7:0] DM_AXI_AWLEN,
    output wire [                 2:0] DM_AXI_AWSIZE,
    output wire [                 1:0] DM_AXI_AWBURST,
    output wire                        DM_AXI_AWLOCK,
    output wire [                 3:0] DM_AXI_AWCACHE,
    output wire [                 2:0] DM_AXI_AWPROT,
    output wire                        DM_AXI_AWVALID,
    input  wire                        DM_AXI_AWREADY,
    output wire [    C_AXI_DATA_WIDTH-1:0] DM_AXI_WDATA,
    output wire [(C_AXI_DATA_WIDTH/8)-1:0] DM_AXI_WSTRB,
    output wire                            DM_AXI_WLAST,
    output wire                            DM_AXI_WVALID,
    input  wire                            DM_AXI_WREADY,
    input  wire [C_AXI_ID_WIDTH-1:0] DM_AXI_BID,
    input  wire [               1:0] DM_AXI_BRESP,
    input  wire                      DM_AXI_BVALID,
    output wire                      DM_AXI_BREADY,
    output wire [  C_AXI_ID_WIDTH-1:0] DM_AXI_ARID,
    output wire [C_AXI_ADDR_WIDTH-1:0] DM_AXI_ARADDR,
    output wire [                 7:0] DM_AXI_ARLEN,
    output wire [                 2:0] DM_AXI_ARSIZE,
    output wire [                 1:0] DM_AXI_ARBURST,
    output wire                        DM_AXI_ARLOCK,
    output wire [                 3:0] DM_AXI_ARCACHE,
    output wire [                 2:0] DM_AXI_ARPROT,
    output wire                        DM_AXI_ARVALID,
    input  wire                        DM_AXI_ARREADY,
    input  wire [  C_AXI_ID_WIDTH-1:0] DM_AXI_RID,
    input  wire [C_AXI_DATA_WIDTH-1:0] DM_AXI_RDATA,
    input  wire [                 1:0] DM_AXI_RRESP,
    input  wire                        DM_AXI_RLAST,
    input  wire                        DM_AXI_RVALID,
    output wire                        DM_AXI_RREADY
);

    // MUX和Crossbar之间的连线
    wire [C_AXI_ID_WIDTH-1:0]     mux_s_axi_awid;
    wire [C_AXI_ADDR_WIDTH-1:0]  mux_s_axi_awaddr;
    wire [7:0]                    mux_s_axi_awlen;
    wire [2:0]                    mux_s_axi_awsize;
    wire [1:0]                    mux_s_axi_awburst;
    wire                          mux_s_axi_awlock;
    wire [3:0]                    mux_s_axi_awcache;
    wire [2:0]                    mux_s_axi_awprot;
    wire [3:0]                    mux_s_axi_awqos;
    wire [3:0]                    mux_s_axi_awuser;
    wire                          mux_s_axi_awvalid;
    wire                          mux_s_axi_awready;
    wire [C_AXI_DATA_WIDTH-1:0]  mux_s_axi_wdata;
    wire [(C_AXI_DATA_WIDTH/8)-1:0] mux_s_axi_wstrb;
    wire                          mux_s_axi_wlast;
    wire                          mux_s_axi_wvalid;
    wire                          mux_s_axi_wready;
    wire [C_AXI_ID_WIDTH-1:0]     mux_s_axi_bid;
    wire [1:0]                    mux_s_axi_bresp;
    wire                          mux_s_axi_bvalid;
    wire                          mux_s_axi_bready;
    wire [C_AXI_ID_WIDTH-1:0]     mux_s_axi_arid;
    wire [C_AXI_ADDR_WIDTH-1:0]  mux_s_axi_araddr;
    wire [7:0]                    mux_s_axi_arlen;
    wire [2:0]                    mux_s_axi_arsize;
    wire [1:0]                    mux_s_axi_arburst;
    wire                          mux_s_axi_arlock;
    wire [3:0]                    mux_s_axi_arcache;
    wire [2:0]                    mux_s_axi_arprot;
    wire [3:0]                    mux_s_axi_arqos;
    wire [3:0]                    mux_s_axi_aruser;
    wire                          mux_s_axi_arvalid;
    wire                          mux_s_axi_arready;
    wire [C_AXI_ID_WIDTH-1:0]     mux_s_axi_rid;
    wire [C_AXI_DATA_WIDTH-1:0]  mux_s_axi_rdata;
    wire [1:0]                    mux_s_axi_rresp;
    wire                          mux_s_axi_rlast;
    wire [3:0]                    mux_s_axi_ruser;
    wire                          mux_s_axi_rvalid;
    wire                          mux_s_axi_rready;

    axi_master_mux #(
        .C_AXI_ID_WIDTH(C_AXI_ID_WIDTH),
        .C_AXI_DATA_WIDTH(C_AXI_DATA_WIDTH),
        .C_AXI_ADDR_WIDTH(C_AXI_ADDR_WIDTH)
    ) i_axi_master_mux (
        .clk(clk),
        .rst_n(rst_n),

        .M0_AXI_ARID(M0_AXI_ARID),
        .M0_AXI_ARADDR(M0_AXI_ARADDR),
        .M0_AXI_ARLEN(M0_AXI_ARLEN),
        .M0_AXI_ARSIZE(M0_AXI_ARSIZE),
        .M0_AXI_ARBURST(M0_AXI_ARBURST),
        .M0_AXI_ARLOCK(M0_AXI_ARLOCK),
        .M0_AXI_ARCACHE(M0_AXI_ARCACHE),
        .M0_AXI_ARPROT(M0_AXI_ARPROT),
        .M0_AXI_ARQOS(M0_AXI_ARQOS),
        .M0_AXI_ARUSER(M0_AXI_ARUSER),
        .M0_AXI_ARVALID(M0_AXI_ARVALID),
        .M0_AXI_ARREADY(M0_AXI_ARREADY),
        .M0_AXI_RID(M0_AXI_RID),
        .M0_AXI_RDATA(M0_AXI_RDATA),
        .M0_AXI_RRESP(M0_AXI_RRESP),
        .M0_AXI_RLAST(M0_AXI_RLAST),
        .M0_AXI_RUSER(M0_AXI_RUSER),
        .M0_AXI_RVALID(M0_AXI_RVALID),
        .M0_AXI_RREADY(M0_AXI_RREADY),

        .M1_AXI_AWID(M1_AXI_AWID),
        .M1_AXI_AWADDR(M1_AXI_AWADDR),
        .M1_AXI_AWLEN(M1_AXI_AWLEN),
        .M1_AXI_AWSIZE(M1_AXI_AWSIZE),
        .M1_AXI_AWBURST(M1_AXI_AWBURST),
        .M1_AXI_AWLOCK(M1_AXI_AWLOCK),
        .M1_AXI_AWCACHE(M1_AXI_AWCACHE),
        .M1_AXI_AWPROT(M1_AXI_AWPROT),
        .M1_AXI_AWQOS(M1_AXI_AWQOS),
        .M1_AXI_AWUSER(M1_AXI_AWUSER),
        .M1_AXI_AWVALID(M1_AXI_AWVALID),
        .M1_AXI_AWREADY(M1_AXI_AWREADY),
        .M1_AXI_WDATA(M1_AXI_WDATA),
        .M1_AXI_WSTRB(M1_AXI_WSTRB),
        .M1_AXI_WLAST(M1_AXI_WLAST),
        .M1_AXI_WVALID(M1_AXI_WVALID),
        .M1_AXI_WREADY(M1_AXI_WREADY),
        .M1_AXI_BID(M1_AXI_BID),
        .M1_AXI_BRESP(M1_AXI_BRESP),
        .M1_AXI_BVALID(M1_AXI_BVALID),
        .M1_AXI_BREADY(M1_AXI_BREADY),
        .M1_AXI_ARID(M1_AXI_ARID),
        .M1_AXI_ARADDR(M1_AXI_ARADDR),
        .M1_AXI_ARLEN(M1_AXI_ARLEN),
        .M1_AXI_ARSIZE(M1_AXI_ARSIZE),
        .M1_AXI_ARBURST(M1_AXI_ARBURST),
        .M1_AXI_ARLOCK(M1_AXI_ARLOCK),
        .M1_AXI_ARCACHE(M1_AXI_ARCACHE),
        .M1_AXI_ARPROT(M1_AXI_ARPROT),
        .M1_AXI_ARQOS(M1_AXI_ARQOS),
        .M1_AXI_ARUSER(M1_AXI_ARUSER),
        .M1_AXI_ARVALID(M1_AXI_ARVALID),
        .M1_AXI_ARREADY(M1_AXI_ARREADY),
        .M1_AXI_RID(M1_AXI_RID),
        .M1_AXI_RDATA(M1_AXI_RDATA),
        .M1_AXI_RRESP(M1_AXI_RRESP),
        .M1_AXI_RLAST(M1_AXI_RLAST),
        .M1_AXI_RUSER(M1_AXI_RUSER),
        .M1_AXI_RVALID(M1_AXI_RVALID),
        .M1_AXI_RREADY(M1_AXI_RREADY),

        .S_AXI_AWID(mux_s_axi_awid),
        .S_AXI_AWADDR(mux_s_axi_awaddr),
        .S_AXI_AWLEN(mux_s_axi_awlen),
        .S_AXI_AWSIZE(mux_s_axi_awsize),
        .S_AXI_AWBURST(mux_s_axi_awburst),
        .S_AXI_AWLOCK(mux_s_axi_awlock),
        .S_AXI_AWCACHE(mux_s_axi_awcache),
        .S_AXI_AWPROT(mux_s_axi_awprot),
        .S_AXI_AWQOS(mux_s_axi_awqos),
        .S_AXI_AWUSER(mux_s_axi_awuser),
        .S_AXI_AWVALID(mux_s_axi_awvalid),
        .S_AXI_AWREADY(mux_s_axi_awready),
        .S_AXI_WDATA(mux_s_axi_wdata),
        .S_AXI_WSTRB(mux_s_axi_wstrb),
        .S_AXI_WLAST(mux_s_axi_wlast),
        .S_AXI_WVALID(mux_s_axi_wvalid),
        .S_AXI_WREADY(mux_s_axi_wready),
        .S_AXI_BID(mux_s_axi_bid),
        .S_AXI_BRESP(mux_s_axi_bresp),
        .S_AXI_BVALID(mux_s_axi_bvalid),
        .S_AXI_BREADY(mux_s_axi_bready),
        .S_AXI_ARID(mux_s_axi_arid),
        .S_AXI_ARADDR(mux_s_axi_araddr),
        .S_AXI_ARLEN(mux_s_axi_arlen),
        .S_AXI_ARSIZE(mux_s_axi_arsize),
        .S_AXI_ARBURST(mux_s_axi_arburst),
        .S_AXI_ARLOCK(mux_s_axi_arlock),
        .S_AXI_ARCACHE(mux_s_axi_arcache),
        .S_AXI_ARPROT(mux_s_axi_arprot),
        .S_AXI_ARQOS(mux_s_axi_arqos),
        .S_AXI_ARUSER(mux_s_axi_aruser),
        .S_AXI_ARVALID(mux_s_axi_arvalid),
        .S_AXI_ARREADY(mux_s_axi_arready),
        .S_AXI_RID(mux_s_axi_rid),
        .S_AXI_RDATA(mux_s_axi_rdata),
        .S_AXI_RRESP(mux_s_axi_rresp),
        .S_AXI_RLAST(mux_s_axi_rlast),
        .S_AXI_RUSER(mux_s_axi_ruser),
        .S_AXI_RVALID(mux_s_axi_rvalid),
        .S_AXI_RREADY(mux_s_axi_rready)
    );

    axi_crossbar #(
        .IMEM_ADDR_WIDTH(IMEM_ADDR_WIDTH),
        .DMEM_ADDR_WIDTH(DMEM_ADDR_WIDTH),
        .DATA_WIDTH(DATA_WIDTH),
        .C_AXI_ID_WIDTH(C_AXI_ID_WIDTH),
        .C_AXI_DATA_WIDTH(C_AXI_DATA_WIDTH),
        .C_AXI_ADDR_WIDTH(C_AXI_ADDR_WIDTH),
        .C_OM0_AXI_ADDR_WIDTH(C_OM0_AXI_ADDR_WIDTH),
        .C_OM0_AXI_DATA_WIDTH(C_OM0_AXI_DATA_WIDTH),
        .C_OM1_AXI_ADDR_WIDTH(C_OM1_AXI_ADDR_WIDTH),
        .C_OM1_AXI_DATA_WIDTH(C_OM1_AXI_DATA_WIDTH),
        .C_OM2_AXI_ADDR_WIDTH(C_OM2_AXI_ADDR_WIDTH),
        .C_OM2_AXI_DATA_WIDTH(C_OM2_AXI_DATA_WIDTH)
    ) i_axi_crossbar (
        .clk(clk),
        .rst_n(rst_n),

        .S_AXI_AWID(mux_s_axi_awid),
        .S_AXI_AWADDR(mux_s_axi_awaddr),
        .S_AXI_AWLEN(mux_s_axi_awlen),
        .S_AXI_AWSIZE(mux_s_axi_awsize),
        .S_AXI_AWBURST(mux_s_axi_awburst),
        .S_AXI_AWLOCK(mux_s_axi_awlock),
        .S_AXI_AWCACHE(mux_s_axi_awcache),
        .S_AXI_AWPROT(mux_s_axi_awprot),
        .S_AXI_AWQOS(mux_s_axi_awqos),
        .S_AXI_AWUSER(mux_s_axi_awuser),
        .S_AXI_AWVALID(mux_s_axi_awvalid),
        .S_AXI_AWREADY(mux_s_axi_awready),
        .S_AXI_WDATA(mux_s_axi_wdata),
        .S_AXI_WSTRB(mux_s_axi_wstrb),
        .S_AXI_WLAST(mux_s_axi_wlast),
        .S_AXI_WVALID(mux_s_axi_wvalid),
        .S_AXI_WREADY(mux_s_axi_wready),
        .S_AXI_BID(mux_s_axi_bid),
        .S_AXI_BRESP(mux_s_axi_bresp),
        .S_AXI_BVALID(mux_s_axi_bvalid),
        .S_AXI_BREADY(mux_s_axi_bready),
        .S_AXI_ARID(mux_s_axi_arid),
        .S_AXI_ARADDR(mux_s_axi_araddr),
        .S_AXI_ARLEN(mux_s_axi_arlen),
        .S_AXI_ARSIZE(mux_s_axi_arsize),
        .S_AXI_ARBURST(mux_s_axi_arburst),
        .S_AXI_ARLOCK(mux_s_axi_arlock),
        .S_AXI_ARCACHE(mux_s_axi_arcache),
        .S_AXI_ARPROT(mux_s_axi_arprot),
        .S_AXI_ARQOS(mux_s_axi_arqos),
        .S_AXI_ARUSER(mux_s_axi_aruser),
        .S_AXI_ARVALID(mux_s_axi_arvalid),
        .S_AXI_ARREADY(mux_s_axi_arready),
        .S_AXI_RID(mux_s_axi_rid),
        .S_AXI_RDATA(mux_s_axi_rdata),
        .S_AXI_RRESP(mux_s_axi_rresp),
        .S_AXI_RLAST(mux_s_axi_rlast),
        .S_AXI_RUSER(mux_s_axi_ruser),
        .S_AXI_RVALID(mux_s_axi_rvalid),
        .S_AXI_RREADY(mux_s_axi_rready),

        .OM0_AXI_ACLK(OM0_AXI_ACLK),
        .OM0_AXI_ARESETN(OM0_AXI_ARESETN),
        .OM0_AXI_AWADDR(OM0_AXI_AWADDR),
        .OM0_AXI_AWPROT(OM0_AXI_AWPROT),
        .OM0_AXI_AWVALID(OM0_AXI_AWVALID),
        .OM0_AXI_AWREADY(OM0_AXI_AWREADY),
        .OM0_AXI_WDATA(OM0_AXI_WDATA),
        .OM0_AXI_WSTRB(OM0_AXI_WSTRB),
        .OM0_AXI_WVALID(OM0_AXI_WVALID),
        .OM0_AXI_WREADY(OM0_AXI_WREADY),
        .OM0_AXI_BRESP(OM0_AXI_BRESP),
        .OM0_AXI_BVALID(OM0_AXI_BVALID),
        .OM0_AXI_BREADY(OM0_AXI_BREADY),
        .OM0_AXI_ARADDR(OM0_AXI_ARADDR),
        .OM0_AXI_ARPROT(OM0_AXI_ARPROT),
        .OM0_AXI_ARVALID(OM0_AXI_ARVALID),
        .OM0_AXI_ARREADY(OM0_AXI_ARREADY),
        .OM0_AXI_RDATA(OM0_AXI_RDATA),
        .OM0_AXI_RRESP(OM0_AXI_RRESP),
        .OM0_AXI_RVALID(OM0_AXI_RVALID),
        .OM0_AXI_RREADY(OM0_AXI_RREADY),
        .OM1_AXI_ACLK(OM1_AXI_ACLK),
        .OM1_AXI_ARESETN(OM1_AXI_ARESETN),
        .OM1_AXI_AWADDR(OM1_AXI_AWADDR),
        .OM1_AXI_AWPROT(OM1_AXI_AWPROT),
        .OM1_AXI_AWVALID(OM1_AXI_AWVALID),
        .OM1_AXI_AWREADY(OM1_AXI_AWREADY),
        .OM1_AXI_WDATA(OM1_AXI_WDATA),
        .OM1_AXI_WSTRB(OM1_AXI_WSTRB),
        .OM1_AXI_WVALID(OM1_AXI_WVALID),
        .OM1_AXI_WREADY(OM1_AXI_WREADY),
        .OM1_AXI_BRESP(OM1_AXI_BRESP),
        .OM1_AXI_BVALID(OM1_AXI_BVALID),
        .OM1_AXI_BREADY(OM1_AXI_BREADY),
        .OM1_AXI_ARADDR(OM1_AXI_ARADDR),
        .OM1_AXI_ARPROT(OM1_AXI_ARPROT),
        .OM1_AXI_ARVALID(OM1_AXI_ARVALID),
        .OM1_AXI_ARREADY(OM1_AXI_ARREADY),
        .OM1_AXI_RDATA(OM1_AXI_RDATA),
        .OM1_AXI_RRESP(OM1_AXI_RRESP),
        .OM1_AXI_RVALID(OM1_AXI_RVALID),
        .OM1_AXI_RREADY(OM1_AXI_RREADY),
        .OM2_AXI_ACLK(OM2_AXI_ACLK),
        .OM2_AXI_ARESETN(OM2_AXI_ARESETN),
        .OM2_AXI_AWADDR(OM2_AXI_AWADDR),
        .OM2_AXI_AWPROT(OM2_AXI_AWPROT),
        .OM2_AXI_AWVALID(OM2_AXI_AWVALID),
        .OM2_AXI_AWREADY(OM2_AXI_AWREADY),
        .OM2_AXI_WDATA(OM2_AXI_WDATA),
        .OM2_AXI_WSTRB(OM2_AXI_WSTRB),
        .OM2_AXI_WVALID(OM2_AXI_WVALID),
        .OM2_AXI_WREADY(OM2_AXI_WREADY),
        .OM2_AXI_BRESP(OM2_AXI_BRESP),
        .OM2_AXI_BVALID(OM2_AXI_BVALID),
        .OM2_AXI_BREADY(OM2_AXI_BREADY),
        .OM2_AXI_ARADDR(OM2_AXI_ARADDR),
        .OM2_AXI_ARPROT(OM2_AXI_ARPROT),
        .OM2_AXI_ARVALID(OM2_AXI_ARVALID),
        .OM2_AXI_ARREADY(OM2_AXI_ARREADY),
        .OM2_AXI_RDATA(OM2_AXI_RDATA),
        .OM2_AXI_RRESP(OM2_AXI_RRESP),
        .OM2_AXI_RVALID(OM2_AXI_RVALID),
        .OM2_AXI_RREADY(OM2_AXI_RREADY),

        .IMEM_AXI_AWID(IMEM_AXI_AWID),
        .IMEM_AXI_AWADDR(IMEM_AXI_AWADDR),
        .IMEM_AXI_AWLEN(IMEM_AXI_AWLEN),
        .IMEM_AXI_AWSIZE(IMEM_AXI_AWSIZE),
        .IMEM_AXI_AWBURST(IMEM_AXI_AWBURST),
        .IMEM_AXI_AWLOCK(IMEM_AXI_AWLOCK),
        .IMEM_AXI_AWCACHE(IMEM_AXI_AWCACHE),
        .IMEM_AXI_AWPROT(IMEM_AXI_AWPROT),
        .IMEM_AXI_AWVALID(IMEM_AXI_AWVALID),
        .IMEM_AXI_AWREADY(IMEM_AXI_AWREADY),
        .IMEM_AXI_WDATA(IMEM_AXI_WDATA),
        .IMEM_AXI_WSTRB(IMEM_AXI_WSTRB),
        .IMEM_AXI_WLAST(IMEM_AXI_WLAST),
        .IMEM_AXI_WVALID(IMEM_AXI_WVALID),
        .IMEM_AXI_WREADY(IMEM_AXI_WREADY),
        .IMEM_AXI_BID(IMEM_AXI_BID),
        .IMEM_AXI_BRESP(IMEM_AXI_BRESP),
        .IMEM_AXI_BVALID(IMEM_AXI_BVALID),
        .IMEM_AXI_BREADY(IMEM_AXI_BREADY),
        .IMEM_AXI_ARID(IMEM_AXI_ARID),
        .IMEM_AXI_ARADDR(IMEM_AXI_ARADDR),
        .IMEM_AXI_ARLEN(IMEM_AXI_ARLEN),
        .IMEM_AXI_ARSIZE(IMEM_AXI_ARSIZE),
        .IMEM_AXI_ARBURST(IMEM_AXI_ARBURST),
        .IMEM_AXI_ARLOCK(IMEM_AXI_ARLOCK),
        .IMEM_AXI_ARCACHE(IMEM_AXI_ARCACHE),
        .IMEM_AXI_ARPROT(IMEM_AXI_ARPROT),
        .IMEM_AXI_ARVALID(IMEM_AXI_ARVALID),
        .IMEM_AXI_ARREADY(IMEM_AXI_ARREADY),
        .IMEM_AXI_RID(IMEM_AXI_RID),
        .IMEM_AXI_RDATA(IMEM_AXI_RDATA),
        .IMEM_AXI_RRESP(IMEM_AXI_RRESP),
        .IMEM_AXI_RLAST(IMEM_AXI_RLAST),
        .IMEM_AXI_RVALID(IMEM_AXI_RVALID),
        .IMEM_AXI_RREADY(IMEM_AXI_RREADY),

        .DMEM_AXI_AWID(DMEM_AXI_AWID),
        .DMEM_AXI_AWADDR(DMEM_AXI_AWADDR),
        .DMEM_AXI_AWLEN(DMEM_AXI_AWLEN),
        .DMEM_AXI_AWSIZE(DMEM_AXI_AWSIZE),
        .DMEM_AXI_AWBURST(DMEM_AXI_AWBURST),
        .DMEM_AXI_AWLOCK(DMEM_AXI_AWLOCK),
        .DMEM_AXI_AWCACHE(DMEM_AXI_AWCACHE),
        .DMEM_AXI_AWPROT(DMEM_AXI_AWPROT),
        .DMEM_AXI_AWVALID(DMEM_AXI_AWVALID),
        .DMEM_AXI_AWREADY(DMEM_AXI_AWREADY),
        .DMEM_AXI_WDATA(DMEM_AXI_WDATA),
        .DMEM_AXI_WSTRB(DMEM_AXI_WSTRB),
        .DMEM_AXI_WLAST(DMEM_AXI_WLAST),
        .DMEM_AXI_WVALID(DMEM_AXI_WVALID),
        .DMEM_AXI_WREADY(DMEM_AXI_WREADY),
        .DMEM_AXI_BID(DMEM_AXI_BID),
        .DMEM_AXI_BRESP(DMEM_AXI_BRESP),
        .DMEM_AXI_BVALID(DMEM_AXI_BVALID),
        .DMEM_AXI_BREADY(DMEM_AXI_BREADY),
        .DMEM_AXI_ARID(DMEM_AXI_ARID),
        .DMEM_AXI_ARADDR(DMEM_AXI_ARADDR),
        .DMEM_AXI_ARLEN(DMEM_AXI_ARLEN),
        .DMEM_AXI_ARSIZE(DMEM_AXI_ARSIZE),
        .DMEM_AXI_ARBURST(DMEM_AXI_ARBURST),
        .DMEM_AXI_ARLOCK(DMEM_AXI_ARLOCK),
        .DMEM_AXI_ARCACHE(DMEM_AXI_ARCACHE),
        .DMEM_AXI_ARPROT(DMEM_AXI_ARPROT),
        .DMEM_AXI_ARVALID(DMEM_AXI_ARVALID),
        .DMEM_AXI_ARREADY(DMEM_AXI_ARREADY),
        .DMEM_AXI_RID(DMEM_AXI_RID),
        .DMEM_AXI_RDATA(DMEM_AXI_RDATA),
        .DMEM_AXI_RRESP(DMEM_AXI_RRESP),
        .DMEM_AXI_RLAST(DMEM_AXI_RLAST),
        .DMEM_AXI_RVALID(DMEM_AXI_RVALID),
        .DMEM_AXI_RREADY(DMEM_AXI_RREADY),

        .DM_AXI_AWID(DM_AXI_AWID),
        .DM_AXI_AWADDR(DM_AXI_AWADDR),
        .DM_AXI_AWLEN(DM_AXI_AWLEN),
        .DM_AXI_AWSIZE(DM_AXI_AWSIZE),
        .DM_AXI_AWBURST(DM_AXI_AWBURST),
        .DM_AXI_AWLOCK(DM_AXI_AWLOCK),
        .DM_AXI_AWCACHE(DM_AXI_AWCACHE),
        .DM_AXI_AWPROT(DM_AXI_AWPROT),
        .DM_AXI_AWVALID(DM_AXI_AWVALID),
        .DM_AXI_AWREADY(DM_AXI_AWREADY),
        .DM_AXI_WDATA(DM_AXI_WDATA),
        .DM_AXI_WSTRB(DM_AXI_WSTRB),
        .DM_AXI_WLAST(DM_AXI_WLAST),
        .DM_AXI_WVALID(DM_AXI_WVALID),
        .DM_AXI_WREADY(DM_AXI_WREADY),
        .DM_AXI_BID(DM_AXI_BID),
        .DM_AXI_BRESP(DM_AXI_BRESP),
        .DM_AXI_BVALID(DM_AXI_BVALID),
        .DM_AXI_BREADY(DM_AXI_BREADY),
        .DM_AXI_ARID(DM_AXI_ARID),
        .DM_AXI_ARADDR(DM_AXI_ARADDR),
        .DM_AXI_ARLEN(DM_AXI_ARLEN),
        .DM_AXI_ARSIZE(DM_AXI_ARSIZE),
        .DM_AXI_ARBURST(DM_AXI_ARBURST),
        .DM_AXI_ARLOCK(DM_AXI_ARLOCK),
        .DM_AXI_ARCACHE(DM_AXI_ARCACHE),
        .DM_AXI_ARPROT(DM_AXI_ARPROT),
        .DM_AXI_ARVALID(DM_AXI_ARVALID),
        .DM_AXI_ARREADY(DM_AXI_ARREADY),
        .DM_AXI_RID(DM_AXI_RID),
        .DM_AXI_RDATA(DM_AXI_RDATA),
        .DM_AXI_RRESP(DM_AXI_RRESP),
        .DM_AXI_RLAST(DM_AXI_RLAST),
        .DM_AXI_RVALID(DM_AXI_RVALID),
        .DM_AXI_RREADY(DM_AXI_RREADY)
    );

endmodule
